----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/03/2024 05:19:30 PM
-- Design Name: 
-- Module Name: ROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;


entity ROM is
    generic
        (
    N_data    : natural := 2;
    N_addr    : natural := 9
        );
    Port ( clk : in STD_LOGIC;
           address : in STD_LOGIC_VECTOR (N_addr-1 downto 0);
           data : out STD_LOGIC_VECTOR (N_data-1 downto 0));
end ROM;

architecture Behavioral of ROM is
  -- type memoire : tableau de 2**N_addr donnees de N_data bits
  type memory_type is array (0 to 2**(N_addr)-1) of std_logic_vector (N_data-1 downto 0); 
  
  
  -- definition du contenu de la memoire
  constant memory_values : memory_type := ("1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","1011","1111","1011","1011","0010","0010","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0000","0010","0000","1000","1111","1010","1111","1010","0000","0000","0000","0000","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","1100","0011","0010","1000","1111","0011","0010","1000","1111","1010","1111","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0000","0000","0000","0000","0011","0010","1100","1000","0011","0010","1100","1000","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0011","1111","0010","1010","0000","0010","0010","0010","1000","0000","0011","1100","1010","1011","0001","1001","1111","0111","0101","0100","1100","1000","0011","0010","1000","1100","1111","1011","1010","0000","1000","1100","0011","1100","1010","1111","1100","1110","1010","0010","1010","1111","1010","1111","1010","1111","1110","0110","0000","1010","0101","0010","1000","1100","1111","1101","1001","1011","1000","1010","1111","0101","1011","1010","0101","0110","1010","1000","1111","0011","1011","1010","1110","1100","1101","0101","0001","0011","0011","0000","0000","1100","0111","0010","0010","1000","1000","1010","1000","1100","1111","1111","0111","0010","1010","1000","1100","1011","1000","1001","0110","0000","0001","1111","1110","0110","0010","0011","1111","1101","1100","1000","1001","1111","0110","1010","0101","0100","1101","0100","1101","0100","1101","0100","1101","1010","0101","1010","0101","1010","0101","1010","0101","0101","1111","1111","1111","1010","1000","1010","1000","1111","1010","1000","1010","1000","1111","1110","1111","1011","1100","1111","1110","1111","1010","1000","1010","1000","1111","1010","1000","1010","1000","1111","1110","1111","1010","1000","1010","1000","1111","1010","1000","1010","1010","1000","1000","1111","1110","1111","1010","1000","1010","1000","1111","1010","1010","1000","1000","1010","1000","1101","1100","1011","1100","1101","1010","1010","1000","1000","1010","1000","1111","1110","1111","1010","1000","1010","1000","1111","1110","1111","1010","1000","1010","1000","1111","1010","1000","1010","1000","1111","1110","1111","1011","1100","1111","1110","1111","1010","1000","1010","1000","1111","1010","1000","1010","1000","1111","1110","1111","1010","1000","1010","1000","1111","1010","1000","1010","1000","1111","1110","1111","1010","1000","1010","1000","1111","1010");
begin  
   -- description ROM synchrone
  process(clk) is
  begin 
    if rising_edge(clk) then      
      data <= memory_values(to_integer(unsigned(address)));           
    end if;
  end process;
end Behavioral;
